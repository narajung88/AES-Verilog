module AES_Generators